
// scoreboard: checks if the cpu is working
class scoreboard;

    

endclass


