// coverage: captures functional coverage information
class coverage;

    virtual cpu_bfm bfm;

endclass
